/********1*********2*********3*********4*********5*********6*********7*********8
*
* FILE      : hex2seg.v
* FUNCTION  : 7-seg display De2-115
* AUTHOR    :
*
*_______________________________________________________________________________
*
* REVISION HISTORY
*
* Name                 Date         Comments
* ------------------------------------------------------------------------------
* oalonso           xx/March/2014     Created
* ------------------------------------------------------------------------------
*_______________________________________________________________________________
* 
* FUNCTIONAL DESCRIPTION 
*
*_______________________________________________________________________________
* 
* (c) Copyright Universitat de Barcelona, 2014 
* All rights reserved. Copying or other reproduction of this 
* program except for archival purposes is prohibited.
*
*********1*********2*********3*********4*********5*********6*********7*********/

module hex2seg(
Clk,Data, Rst_n, seg
);
input Clk, Rst_n;
output [7:0] seg;
input [3:0] Data;
reg [7:0] seg;


always @(posedge Clk or negedge Rst_n)
	case(Data)
		4'd0: seg[7:0] <= ~(8'b00111111);
		4'd1: seg[7:0] <= ~(8'b00000110);
		4'd2: seg[7:0] <= ~(8'b01011011);
		4'd3: seg[7:0] <= ~(8'b01001111);
		4'd4: seg[7:0] <= ~(8'b01100110);
		4'd5: seg[7:0] <= ~(8'b01101101);
		4'd6: seg[7:0] <= ~(8'b01111101);
		4'd7: seg[7:0] <= ~(8'b00000111);
		4'd8: seg[7:0] <= ~(8'b01111111);
		4'd9: seg[7:0] <= ~(8'b01100111);
		4'hA: seg[7:0] <= ~(8'b01110111);
		4'hB: seg[7:0] <= ~(8'b01111100);
		4'hC: seg[7:0] <= ~(8'b00111001);
		4'hD: seg[7:0] <= ~(8'b01011110);
		4'hE: seg[7:0] <= ~(8'b01111001);
		4'hF: seg[7:0] <= ~(8'b01110001);
	endcase

endmodule
